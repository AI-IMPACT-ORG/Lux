Require Import M3Coq RGCoq TestsCoq MultiLogicBundle Metalogic.

(* Aggregate module for convenience. *)
